
module matrix_mul (
	clk_clk);	

	input		clk_clk;
endmodule
