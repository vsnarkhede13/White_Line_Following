
module hello_world (
	clk_clk);	

	input		clk_clk;
endmodule
